module Controler (opcode,func,clock,Reset,PCWrite,IorD,MemWrite,MemToReg,IRWrite,PCSrc,ALUop,ALUSrcA,ALUSrcB,RegWrite,RegDst,ALUout,AWrite,BWrite);
	input wire [5:0] opcode,func;
	input wire clock;
	reg [5:0] Fetch,Wait1,InstRead,Wait2,OpcodeRead,WriteRegALU,ResetS;
	output reg Reset,PCWrite,MemWrite,IRWrite,RegWrite,ALUout,AWrite,BWrite;
	output reg [1:0] ALUSrcA,RegDst;
	output reg [2:0] IorD,PCSrc,ALUop,ALUSrcB;
	output reg [3:0] MemToReg;
	reg [5:0] Estado;
	initial begin 
		Estado <= 6'd0;
		ResetS <= 6'd0;
		Fetch <= 6'd1;
		Wait1 <= 6'd2;
		InstRead <= 6'd3;
		Wait2 <= 6'd4;
		OpcodeRead <= 6'd5;
		WriteRegALU <= 6'd6;
	end
	
		
	always @(posedge clock) begin
		case(Estado)
			ResetS: begin
				Reset <= 1'b1;
				Estado <= Fetch;
			end
			Fetch: begin //Solicita Leitura da Memoria e faz PC + 4
				PCWrite <= 1'b1;
				PCSrc <= 3'b000;
				ALUop <= 3'b001;
				ALUSrcA <= 2'b00;
				AWrite <= 1'b1;
				ALUSrcB <= 3'b001;
				BWrite <= 1'b1;
				Reset <= 1'b0;
				IorD <= 3'b100;
				IRWrite <= 1'b0;
				MemWrite <= 1'b0;
				MemToReg <= 4'b0000;
				RegWrite <= 1'b0;
				RegDst <= 2'b00;
				ALUout <= 1'b1;
				Estado <= Wait1;				
			end
			Wait1: begin
				PCWrite <= 1'b0;
				ALUout <= 1'b0;
				AWrite <= 1'b0;
				BWrite <= 1'b0;
				Estado <= InstRead;
			end
			InstRead: begin //Carrega Dados da Memoria nos Registradores de Instru��o e Opera��o (A e B).
				PCWrite <= 1'b0;
				IRWrite <= 1'b1;
				Estado <= Wait2;
			end
			Wait2: begin
				IRWrite <= 1'b0;
				PCWrite <= 1'b0;
				Estado <= OpcodeRead;			
			end
			WriteRegALU: begin
				MemToReg <= 4'b0000;
				RegDst <= 2'b11;
				RegWrite <= 1'b1;
				Estado <= Fetch;
			end
			OpcodeRead: begin
				case(opcode)
					6'd0: begin
						case(func)
							6'b100000: begin //Add
								ALUop <= 3'b001;
								ALUSrcA <= 2'b10;
								ALUSrcB <= 3'b000;
								ALUout <= 1'b1;
								Estado <= WriteRegALU;
							end
						endcase
					end		
				endcase
			end
				
		endcase
	end
endmodule 	